`timescale 1ns / 1ps

module TopModule_Switch
#(
	parameter WIDTH = 128, // larghezza del bundled data.=256
	parameter PORTS =5,
	parameter int BUFNumber [PORTS-1:0]= {6,6,5,7,5},
	parameter int BUFNumberIO [PORTS-1:0]= {4,2,3,4,4}
  
)
(
	input 							 reset,
	input 							 gen_enable,
	
	input			[PORTS-1:0]	req_up_i,
	input			[WIDTH-1:0] Data_up_i_0,
	input			[WIDTH-1:0] Data_up_i_1,
	input			[WIDTH-1:0] Data_up_i_2,
	input			[WIDTH-1:0] Data_up_i_3,
	input			[WIDTH-1:0] Data_up_i_4,
	output		[PORTS-1:0]	ack_up_o,

	output   [PORTS-1:0]req_dw_o,
	output   [WIDTH-1:0] Data_dw0_o,
	output   [WIDTH-1:0] Data_dw1_o,
	output   [WIDTH-1:0] Data_dw2_o,
	output   [WIDTH-1:0] Data_dw3_o,
	output   [WIDTH-1:0] Data_dw4_o,
	input    [PORTS-1:0] ack_dw_i
);

    logic [PORTS-1:0][WIDTH-1:0]  DataAuxIn,DataAuxOut;
    assign DataAuxIn = {Data_up_i_4,Data_up_i_3,Data_up_i_2,Data_up_i_1,Data_up_i_0}; 
    assign DataAuxOut = {Data_dw4_o,Data_dw3_o,Data_dw2_o,Data_dw1_o,Data_dw0_o}; 
    /*
    (* DONT_TOUCH = "yes"*) opm#(WIDTH,PORTS) Myopm(reset,gen_enable,req_up_i,DataAusiliary,ack_up_o,req_dw_o,Data_dw0_o,ack_dw_i,PacketEnable_up_i,Tailpassed_dw_i);
    */
    Switch#(WIDTH,2,2,4,1,BUFNumber,BUFNumberIO) mySwitch(reset,gen_enable,req_up_i,DataAuxIn,ack_up_o,req_dw_o,DataAuxOut,ack_dw_i);
endmodule









































































































































































































































































































































































































































































































































































































































































































































































































































































